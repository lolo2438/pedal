library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity dsp is
end entity;

architecture rtl of dsp is
begin

end architecture;
