library ieee;
use ieee.std_logic_1164.all;

package types_pkg is

  type std_logic_array is array (natural range <>) of std_logic_vector;

end package;
